class dp_seq_a extends uvm_sequencer#(dp_sequence_item_a);
    `uvm_component_utils(dp_seq_a)

    function new(string name = "dp_seq_a",uvm_component parent);
        super.new(name,parent);
    endfunction 

endclass 


